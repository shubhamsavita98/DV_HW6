//`default_nettype none
module my_mem_top(my_mem_inf top_inf);

	my_mem design(top_inf.my_mem);

endmodule